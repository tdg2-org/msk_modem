
package mf_taps_pkg;

  localparam int  MF_NTAPS = 41;

  // 16‑bit half‑sine taps, peak = 32767
  localparam logic signed [15:0] MF_COEFFS [MF_NTAPS] = '{
    16'sd0,      16'sd2571, 16'sd5126, 16'sd7649, 16'sd10126,
    16'sd12539,  16'sd14876, 16'sd17121, 16'sd19260, 16'sd21280,
    16'sd23170,  16'sd24916, 16'sd26509, 16'sd27938, 16'sd29196,
    16'sd30273,  16'sd31163, 16'sd31862, 16'sd32364, 16'sd32666,
    16'sd32767,  16'sd32666, 16'sd32364, 16'sd31862, 16'sd31163,
    16'sd30273,  16'sd29196, 16'sd27938, 16'sd26509, 16'sd24916,
    16'sd23170,  16'sd21280, 16'sd19260, 16'sd17121, 16'sd14876,
    16'sd12539,  16'sd10126, 16'sd7649,  16'sd5126,  16'sd2571,
    16'sd0
  };

endpackage

/* 16bit signed dec

0,2571,5126,7649,10126,12539,14876,17121,19260,21280,23170,24916,26509,27938,29196,30273,31163,31862,32364,32666,32767,32666,32364,31862,31163,30273,29196,27938,26509,24916,23170,21280,19260,17121,14876,12539,10126,7649,5126,2571,0

*/