`timescale 1ns / 1ps  // <time_unit>/<time_precision>

module cfo_test #(
  parameter int SEL = 0,
  parameter int OW  = 16  
)(
  input   logic clk,
  input   logic rst,
  input   logic val,
  output  logic signed [OW-1:0]   i_o,   
  output  logic signed [OW-1:0]   q_o    
);
//-------------------------------------------------------------------------------------------------
// 
//-------------------------------------------------------------------------------------------------
  int sel_i = SEL;

  logic signed [OW-1:0] i0, i1, i2, i3;
  logic signed [OW-1:0] q0, q1, q2, q3;

  assign i_o =  (sel_i == 0) ? i0 :
                (sel_i == 1) ? i1 :
                (sel_i == 2) ? i2 :
                (sel_i == 3) ? i3 :
                '0;

  assign q_o =  (sel_i == 0) ? q0 :
                (sel_i == 1) ? q1 :
                (sel_i == 2) ? q2 :
                (sel_i == 3) ? q3 :
                '0;

//-------------------------------------------------------------------------------------------------
// 
//-------------------------------------------------------------------------------------------------

  int cnt = 0;

  always_ff @(posedge clk) begin
    if (rst) begin 
      //i_sym <= '0;
      //q_sym <= '0;
    end else if (val) begin
      if (cnt == 7) cnt <= '0;
      else cnt <= cnt + 1;
    end 
  end

//-------------------------------------------------------------------------------------------------
// I,Q = (0x7FFF,0) -> (0,0x7FFF) -> (0x8000,0) -> (0,0x8000)
//        (32767,0)     (0,32767)      -32768,0     0,-32768         
// expect freq_word = 0
//-------------------------------------------------------------------------------------------------
  assign i0 = ((cnt == 0) || (cnt == 4)) ? 'h7FFF :
              ((cnt == 1) || (cnt == 5)) ? 0      :
              ((cnt == 2) || (cnt == 6)) ? 'h8000 :
              ((cnt == 3) || (cnt == 7)) ? 0      : 0;
  assign q0 = ((cnt == 0) || (cnt == 4)) ? 0      :
              ((cnt == 1) || (cnt == 5)) ? 'h7FFF :
              ((cnt == 2) || (cnt == 6)) ? 0      :
              ((cnt == 3) || (cnt == 7)) ? 'h8000 : 0;

//-------------------------------------------------------------------------------------------------
// I,Q = (0x7FFF, 0) repeated
//        (32767,0)
// expect freq_word = 0
//-------------------------------------------------------------------------------------------------
  assign i1 = 'h7FFF;
  assign q1 = 0;

//-------------------------------------------------------------------------------------------------
// (0x7FFF,0) (0x5A82,0x5A82) (0,0x7FFF) (‑0x5A82,0x5A82) (-0x7FFF,0x0000) (-0x5A82,-0x5A82) (0x0000,-0x7FFF) (0x5A82,-0x5A82)
// (32767,0)  (23170, 23170)  (0,32767)  (-23170, 23170)
// expect freq_word = 0x2000_0000
//-------------------------------------------------------------------------------------------------
  assign i2 = (cnt == 0) ? 32767  :                     
              (cnt == 1) ? 23170  :                     
              (cnt == 2) ? 0      :                       
              (cnt == 3) ? -23170 :                     
              (cnt == 4) ? -32767 :                          
              (cnt == 5) ? -23170 :                          
              (cnt == 6) ? 0      :                            
              (cnt == 7) ? 23170  : 0;                      

  assign q2 = (cnt == 0) ? 0      :
              (cnt == 1) ? 23170  :
              (cnt == 2) ? 32767  :
              (cnt == 3) ? 23170  :
              (cnt == 4) ? 0      :      
              (cnt == 5) ? -23170 :                
              (cnt == 6) ? -32767 :                
              (cnt == 7) ? -23170 : 0;

  // negate Q, expect freq_word = 0xE000_0000
  assign i3 = (cnt == 0) ? 32767  :                     
              (cnt == 1) ? 23170  :                     
              (cnt == 2) ? 0      :                       
              (cnt == 3) ? -23170 :                     
              (cnt == 4) ? -32767 :                          
              (cnt == 5) ? -23170 :                          
              (cnt == 6) ? 0      :                            
              (cnt == 7) ? 23170  : 0;                      

  assign q3 = (cnt == 0) ? 0      :
              (cnt == 1) ? -23170 :
              (cnt == 2) ? -32767 :
              (cnt == 3) ? -23170 :
              (cnt == 4) ? 0      :      
              (cnt == 5) ? 23170  :                
              (cnt == 6) ? 32767  :                
              (cnt == 7) ? 23170  : 0;


endmodule
/*

  cfo_test #(
    .SEL (0 ),
    .OW  (16)  
  )(
    .clk  (),
    .rst  (),
    .val  (),
    .i_o  (),   
    .q_o  ()    
  );


*/