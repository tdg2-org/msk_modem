
package mf_taps_pkg;

  localparam int MF_NTAPS = 121;

  localparam logic signed [15:0] mf_coeffs [MF_NTAPS-1:0] = {
    -16'd275	,				     
    -16'd232	,				     
    -16'd177	,				     
    -16'd112	,				     
    -16'd37		,			     
    16'd44		,			     
    16'd131		,			     
    16'd221		,			     
    16'd311		,			     
    16'd397		,			     
    16'd478		,			     
    16'd550		,			     
    16'd610		,			     
    16'd655		,			     
    16'd682		,			     
    16'd690		,			     
    16'd676		,			     
    16'd639		,			     
    16'd579		,			     
    16'd495		,			     
    16'd389		,			     
    16'd261		,			     
    16'd115		,			     
    -16'd46		,			     
    -16'd221	,				     
    -16'd403	,				     
    -16'd588	,				     
    -16'd771	,				     
    -16'd946	,				     
    -16'd1107	,				     
    -16'd1249	,				     
    -16'd1364	,				     
    -16'd1447	,				     
    -16'd1494	,				     
    -16'd1499	,				     
    -16'd1457	,				     
    -16'd1366	,				     
    -16'd1223	,				     
    -16'd1026	,				     
    -16'd775	,				     
    -16'd471	,				     
    -16'd115	,				     
    16'd288		,			     
    16'd737		,			     
    16'd1224	,				     
    16'd1744	,				     
    16'd2290	,				     
    16'd2853	,				     
    16'd3425	,				     
    16'd3997	,				     
    16'd4560	,				     
    16'd5105	,				     
    16'd5621	,				     
    16'd6101	,				     
    16'd6536	,				     
    16'd6917	,				     
    16'd7240	,				     
    16'd7497	,				     
    16'd7684	,				     
    16'd7797	,				     
    16'd7835	,				     
    16'd7797	,				     
    16'd7684	,				     
    16'd7497	,				     
    16'd7240	,				     
    16'd6917	,				     
    16'd6536	,				     
    16'd6101	,				     
    16'd5621	,				     
    16'd5105	,				     
    16'd4560	,				     
    16'd3997	,				     
    16'd3425	,				     
    16'd2853	,				     
    16'd2290	,				     
    16'd1744	,				     
    16'd1224	,				     
    16'd737		,			     
    16'd288		,			     
    -16'd115	,				     
    -16'd471	,				     
    -16'd775	,				     
    -16'd1026	,				     
    -16'd1223	,				     
    -16'd1366	,				     
    -16'd1457	,				     
    -16'd1499	,				     
    -16'd1494	,				     
    -16'd1447	,				     
    -16'd1364	,				     
    -16'd1249	,				     
    -16'd1107	,				     
    -16'd946	,				     
    -16'd771	,				     
    -16'd588	,				     
    -16'd403	,				     
    -16'd221	,				     
    -16'd46		,			     
    16'd115		,			     
    16'd261		,			     
    16'd389		,			     
    16'd495		,			     
    16'd579		,			     
    16'd639		,			     
    16'd676		,			     
    16'd690		,			     
    16'd682		,			     
    16'd655		,			     
    16'd610		,			     
    16'd550		,			     
    16'd478		,			     
    16'd397		,			     
    16'd311		,			     
    16'd221		,			     
    16'd131		,			     
    16'd44		,			     
    -16'd37		,			     
    -16'd112	,				     
    -16'd177	,				     
    -16'd232	,				     
    -16'd275	
  };


endpackage
/*
feed		
ff18		
ff4f		
ff90		
ffdb		
002c		
0083		
00dd		
0137		
018d		
01de		
0226		
0262		
028f		
02aa		
02b2		
02a4		
027f		
0243		
01ef		
0185		
0105		
0073		
ffd2		
ff23		
fe6d		
fdb4		
fcfd		
fc4e		
fbad		
fb1f		
faac		
fa59		
fa2a		
fa25		
fa4f		
faaa		
fb39		
fbfe		
fcf9		
fe29		
ff8d		
0120		
02e1		
04c8		
06d0		
08f2		
0b25		
0d61		
0f9d		
11d0		
13f1		
15f5		
17d5		
1988		
1b05		
1c48		
1d49		
1e04		
1e75		
1e9b		
1e75		
1e04		
1d49		
1c48		
1b05		
1988		
17d5		
15f5		
13f1		
11d0		
0f9d		
0d61		
0b25		
08f2		
06d0		
04c8		
02e1		
0120		
ff8d		
fe29		
fcf9		
fbfe		
fb39		
faaa		
fa4f		
fa25		
fa2a		
fa59		
faac		
fb1f		
fbad		
fc4e		
fcfd		
fdb4		
fe6d		
ff23		
ffd2		
0073		
0105		
0185		
01ef		
0243		
027f		
02a4		
02b2		
02aa		
028f		
0262		
0226		
01de		
018d		
0137		
00dd		
0083		
002c		
ffdb		
ff90		
ff4f		
ff18		
feed		
*/


/*BAD:

-16'sd275,
-16'sd232,
-16'sd177,
-16'sd112,
-16'sd38,
16'sd44,
16'sd131,
16'sd221,
16'sd311,
16'sd398,
16'sd479,
16'sd551,
16'sd611,
16'sd655,
16'sd683,
16'sd690,
16'sd677,
16'sd642,
16'sd588,
16'sd515,
16'sd428,
16'sd329,
16'sd221,
16'sd109,
16'sd0,
-16'sd102,
-16'sd195,
-16'sd275,
-16'sd342,
-16'sd392,
-16'sd426,
-16'sd441,
-16'sd438,
-16'sd416,
-16'sd376,
-16'sd318,
-16'sd246,
-16'sd162,
-16'sd70,
16'sd24,
16'sd115,
16'sd201,
16'sd278,
16'sd344,
16'sd397,
16'sd435,
16'sd456,
16'sd461,
16'sd449,
16'sd420,
16'sd377,
16'sd321,
16'sd255,
16'sd184,
16'sd109,
16'sd36,
-16'sd35,
-16'sd99,
-16'sd153,
-16'sd195,
-16'sd222,
-16'sd235,
-16'sd233,
-16'sd217,
-16'sd188,
-16'sd148,
-16'sd99,
-16'sd43,
16'sd14,
16'sd70,
16'sd124,
16'sd170,
16'sd208,
16'sd236,
16'sd252,
16'sd257,
16'sd249,
16'sd229,
16'sd199,
16'sd159,
16'sd111,
16'sd57,
16'sd0,
-16'sd57,
-16'sd111,
-16'sd159,
-16'sd199,
-16'sd229,
-16'sd249,
-16'sd257,
-16'sd252,
-16'sd236,
-16'sd208,
-16'sd170,
-16'sd124,
-16'sd70,
-16'sd14,
16'sd43,
16'sd99,
16'sd148,
16'sd188,
16'sd217,
16'sd233,
16'sd235,
16'sd222,
16'sd195,
16'sd153,
16'sd99,
16'sd35,
-16'sd36,
-16'sd109,
-16'sd184,
-16'sd255,
-16'sd321,
-16'sd377,
-16'sd420,
-16'sd449,
-16'sd461,
-16'sd456,
-16'sd435,
-16'sd397,
-16'sd344,
-16'sd278,
-16'sd201,
-16'sd115,
-16'sd24,
16'sd70,
16'sd162,
16'sd246,
16'sd318,
16'sd376,
16'sd416,
16'sd438,
16'sd441,
16'sd426,
16'sd392,
16'sd342,
16'sd275,
16'sd195,
16'sd102,
16'sd0,
-16'sd109,
-16'sd221,
-16'sd329,
-16'sd428,
-16'sd515,
-16'sd588,
-16'sd642,
-16'sd677,
-16'sd690,
-16'sd683,
-16'sd655,
-16'sd611,
-16'sd551,
-16'sd479,
-16'sd398,
-16'sd311,
-16'sd221,
-16'sd131,
-16'sd44,
16'sd38,
16'sd112,
16'sd177,
16'sd232,
16'sd275

*/
